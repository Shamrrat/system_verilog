modu;uniuic
