module asssertioon;
